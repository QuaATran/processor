//decoder module

module registerDecoder (Dout, selector, enable);

 input enable;					 
 input  [4:0] selector;
 output reg [31:0] Dout;
		  
 always @(posedge enable or posedge selector) begin
  case({selector})
		5'b00000: Dout = 32'b00000000000000000000000000000001;
		5'b00001: Dout = 32'b00000000000000000000000000000010;
		5'b00010: Dout = 32'b00000000000000000000000000000100;
		5'b00011: Dout = 32'b00000000000000000000000000001000;
		5'b00100: Dout = 32'b00000000000000000000000000010000;
		5'b00101: Dout = 32'b00000000000000000000000000100000;
		5'b00110: Dout = 32'b00000000000000000000000001000000;
		5'b00111: Dout = 32'b00000000000000000000000010000000;
		5'b01000: Dout = 32'b00000000000000000000000100000000;
		5'b01001: Dout = 32'b00000000000000000000001000000000;
		5'b01010: Dout = 32'b00000000000000000000010000000000;
		5'b01011: Dout = 32'b00000000000000000000100000000000;
		5'b01100: Dout = 32'b00000000000000000001000000000000;
		5'b01101: Dout = 32'b00000000000000000010000000000000;
		5'b01110: Dout = 32'b00000000000000000100000000000000;
		5'b01111: Dout = 32'b00000000000000001000000000000000;
		5'b10000: Dout = 32'b00000000000000010000000000000000;
		5'b10001: Dout = 32'b00000000000000100000000000000000;
		5'b10010: Dout = 32'b00000000000001000000000000000000;
		5'b10011: Dout = 32'b00000000000010000000000000000000;
		5'b10100: Dout = 32'b00000000000100000000000000000000;
		5'b10101: Dout = 32'b00000000001000000000000000000000;
		5'b10110: Dout = 32'b00000000010000000000000000000000;
		5'b10111: Dout = 32'b00000000100000000000000000000000;
		5'b11000: Dout = 32'b00000001000000000000000000000000;
		5'b11001: Dout = 32'b00000010000000000000000000000000;
		5'b11010: Dout = 32'b00000100000000000000000000000000;
		5'b11011: Dout = 32'b00001000000000000000000000000000;
		5'b11100: Dout = 32'b00010000000000000000000000000000;
		5'b11101: Dout = 32'b00100000000000000000000000000000;
		5'b11110: Dout = 32'b01000000000000000000000000000000;
		5'b11111: Dout = 32'b10000000000000000000000000000000;
	  default: Dout = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
	 endcase
	
	end
	
endmodule 